module ysyx_23060059_clint(
    input   wire         clock,
    input   wire         reset,
    output  wire  [63:0] mtime  
);

    


endmodule